//Your own small assembly-like language +VM for it (+make game with it)

//ref: http://www.ittybittycomputers.com/IttyBitty/IBSM.htm

`ifndef P07__SV

`define P07__SV

 

program P_07;

 

endprogram

 

`endif //P07__SV
